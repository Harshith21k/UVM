module tb;
  int a;
  int b;
  
endmodule
