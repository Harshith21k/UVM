module tb;
  
  
endmodule
